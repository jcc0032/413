module ALU1(In1,In2, Control, theResult);
input [7:0] In1, In2;
input[3:0] Control;
output [7:0] theResult;
// Insert your code here
endmodule